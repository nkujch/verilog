library verilog;
use verilog.vl_types.all;
entity uart_tx_tb is
end uart_tx_tb;
