library verilog;
use verilog.vl_types.all;
entity sys_pll_tb_1 is
end sys_pll_tb_1;
