library verilog;
use verilog.vl_types.all;
entity pll_0_tb is
end pll_0_tb;
